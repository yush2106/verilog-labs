module decoder3to8(
  input wire[2:0] d,
  output wire[7:0] y
);

assign
  y[0] = ~( ~d[2] & ~d[1] & ~d[0] ),    //d[2:0] = 3'b000
  y[1] = ~( ~d[2] & ~d[1] &  d[0] ),    //d[2:0] = 3'b001
  y[2] = ~( ~d[2] &  d[1] & ~d[0] ),    //d[2:0] = 3'b010
  y[3] = ~( ~d[2] &  d[1] &  d[0] ),    //d[2:0] = 3'b011
  y[4] = ~(  d[2] & ~d[1] & ~d[0] ),    //d[2:0] = 3'b100
  y[5] = ~(  d[2] & ~d[1] &  d[0] ),    //d[2:0] = 3'b101
  y[6] = ~(  d[2] &  d[1] & ~d[0] ),    //d[2:0] = 3'b110
  y[7] = ~(  d[2] &  d[1] &  d[0] );    //d[2:0] = 3'b111

endmodule